`define CHAR_WIDTH 8
`define DATA_WIDTH 16

`define QUERY_LEN 101
`define REF_MAX_LEN  1024


